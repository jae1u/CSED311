module ALU #(parameter data_width = 16)
            (input [data_width - 1 : 0] A,
             input [data_width - 1 : 0] B,
             input [3 : 0] FuncCode,
             output reg [data_width - 1: 0] C,
             output reg OverflowFlag);
    // Do not use delay in your implementation.
    
    // You can declare any variables as needed.
    /*
     YOUR VARIABLE DECLARATION...
     */
    
    initial begin
        C            = 0;
        OverflowFlag = 0;
    end
    
    // TODO: You should implement the functionality of ALU!
    // (HINT: Use 'always @(...) begin ... end')
    /*
     YOUR ALU FUNCTIONALITY IMPLEMENTATION...
     */
    
endmodule