`include "def_opcode.v"

module cpu (
    input reset,
    input clk,
    output is_halted,
    output reg [31:0] print_reg [0:31]
);
    /***** Register declarations *****/
    reg [31:0] IR; // instruction register
    reg [31:0] MDR; // memory data register
    reg [31:0] A; // Read 1 data register
    reg [31:0] B; // Read 2 data register
    reg [31:0] ALUOut; // ALU output register
    // Do not modify and use registers declared above.

    // control signals
    wire pc_write;
    wire pc_write_not_cond;
    wire i_or_d;
    wire mem_read;
    wire mem_write;
    wire ir_write;
    wire mem_to_reg;
    wire reg_write;
    wire alu_src_a;
    wire [1:0] alu_src_b;
    wire [1:0] alu_op;
    wire pc_src;
    wire alu_out_write;

    // inter-module wires
    wire pc_actual_write;
    wire [31:0] next_pc;
    wire [31:0] pc_val /* verilator public */;
    wire [31:0] alu_out_val;
    wire [31:0] mem_addr;
    wire [31:0] mem_read_data;
    wire [31:0] ir_val;
    wire [31:0] mdr_val;
    wire [31:0] rf_write_data;
    wire [31:0] rf_read_data_1;
    wire [31:0] rf_read_data_2;
    wire [31:0] read_data_a_val;
    wire [31:0] read_data_b_val;
    wire [31:0] imm;
    wire [3:0] alu_ctl;
    wire [31:0] alu_operand_a;
    wire [31:0] alu_operand_b;
    wire [31:0] alu_result;
    wire bcond;
    wire [31:0] x17_val;
    
    assign pc_actual_write = pc_write | (pc_write_not_cond & ~bcond);
    assign bcond = alu_result[0];
    assign is_halted = (ir_val[6:0] == `ECALL) && (x17_val == 10);

    d_reg pc(
        .reset(reset),
        .data(next_pc),
        .write(pc_actual_write),
        .clk(clk),
        .out(pc_val)
    );

    mux #(.K(32)) mem_addr_mux(
        .ins({alu_out_val, pc_val}),
        .select(i_or_d),
        .out(mem_addr)
    );

    Memory memory_mod(
        .reset(reset),
        .clk(clk),
        .addr(mem_addr),
        .din(read_data_b_val),
        .mem_read(mem_read),
        .mem_write(mem_write),
        .dout(mem_read_data)
    );

    mux #(.K(32)) rf_write_data_mux(
        .ins({mdr_val, alu_out_val}),
        .select(mem_to_reg),
        .out(rf_write_data)
    );

    RegisterFile rf_mod(
        .reset(reset),
        .clk(clk),
        .rs1(ir_val[19:15]),
        .rs2(ir_val[24:20]),
        .rd(ir_val[11:7]),
        .rd_din(rf_write_data),
        .write_enable(reg_write),
        .rs1_dout(rf_read_data_1),
        .rs2_dout(rf_read_data_2),
        .x17(x17_val),
        .print_reg(print_reg)
    );

    imm_gen imm_gen_mod(
        .instr(ir_val),
        .imm(imm)
    );

    alu_control alu_control_mod(
        .alu_op(alu_op),
        .funct({ir_val[30], ir_val[14:12]}),
        .alu_ctl(alu_ctl)
    );

    mux #(.K(32)) alu_operand_a_mux(
        .ins({read_data_a_val, pc_val}),
        .select(alu_src_a),
        .out(alu_operand_a)
    );

    mux #(.N(2), .K(32)) alu_operand_b_mux(
        .ins({0, imm, 4, read_data_b_val}),
        .select(alu_src_b),
        .out(alu_operand_b)
    );

    alu alu_mod(
        .a(alu_operand_a),
        .b(alu_operand_b),
        .alu_ctl(alu_ctl),
        .result(alu_result)
    );

    mux #(.K(32)) next_pc_mux(
        .ins({alu_out_val, alu_result}),
        .select(pc_src),
        .out(next_pc)
    );

    ucontroller ucontroller_mod(
        .opcode(ir_val[6:0]),
        .bcond(bcond),
        .reset(reset),
        .clk(clk),
        .pc_write(pc_write),
        .pc_write_not_cond(pc_write_not_cond),
        .i_or_d(i_or_d),
        .mem_read(mem_read),
        .mem_write(mem_write),
        .ir_write(ir_write),
        .mem_to_reg(mem_to_reg),
        .reg_write(reg_write),
        .alu_src_a(alu_src_a),
        .alu_src_b(alu_src_b),
        .alu_op(alu_op),
        .pc_src(pc_src),
        .alu_out_write(alu_out_write)
    );

    assign ir_val = IR;
    assign mdr_val = MDR;
    assign read_data_a_val = A;
    assign read_data_b_val = B;
    assign alu_out_val = ALUOut;

    always @(posedge clk) begin
        if (reset) begin
            IR <= 0;
            MDR <= 0;
            A <= 0;
            B <= 0;
            ALUOut <= 0;
        end
        else begin
            if (ir_write) IR <= mem_read_data;
            MDR <= mem_read_data;
            A <= rf_read_data_1;
            B <= rf_read_data_2;
            if (alu_out_write) ALUOut <= alu_result;
        end
    end
endmodule
